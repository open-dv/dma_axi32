`include "dma_axi32_defines.v"
`include "dma_axi32_reg_params.v"
`include "dma_axi32_ch_reg_params.v"
`include "dma_axi32_wrap.v"
`include "axi_slave/axi_slave.v"
`include "axi_slave/axi_slave_addr_gen.v"
`include "axi_slave/axi_slave_busy.v"
`include "axi_slave/axi_slave_cmd_fifo.v"
`include "axi_slave/axi_slave_mem.v"
`include "axi_slave/axi_slave_ram.v"
`include "axi_slave/axi_slave_rd_buff.v"
`include "axi_slave/axi_slave_wresp_fifo.v"
`include "axi_slave/prgen_fifo_stub.v"
`include "axi_slave/prgen_rand.v"
`include "dma_axi32.v"
`include "dma_axi32_dual_core.v"
`include "dma_axi32_apb_mux.v"
`include "dma_axi32_reg.v"
`include "dma_axi32_reg_core0.v"
`include "prgen_scatter8_1.v"
`include "dma_axi32_core0_top.v"
`include "dma_axi32_core0.v"
`include "dma_axi32_core0_wdt.v"
`include "dma_axi32_core0_arbiter.v"
`include "dma_axi32_core0_ctrl.v"
`include "dma_axi32_core0_axim_wr.v"
`include "dma_axi32_core0_axim_cmd.v"
`include "dma_axi32_core0_axim_timeout.v"
`include "dma_axi32_core0_axim_wdata.v"
`include "prgen_joint_stall.v"
`include "prgen_fifo.v"
`include "prgen_stall.v"
`include "dma_axi32_core0_axim_resp.v"
`include "dma_axi32_core0_axim_rd.v"
`include "dma_axi32_core0_axim_rdata.v"
`include "dma_axi32_core0_channels.v"
`include "dma_axi32_core0_channels_apb_mux.v"
`include "dma_axi32_core0_channels_mux.v"
`include "prgen_or8.v"
`include "prgen_mux8.v"
`include "prgen_demux8.v"
`include "dma_axi32_core0_ch.v"
`include "dma_axi32_core0_ch_reg.v"
`include "dma_axi32_core0_ch_reg_size.v"
`include "prgen_rawstat.v"
`include "dma_axi32_core0_ch_offsets.v"
`include "dma_axi32_core0_ch_remain.v"
`include "dma_axi32_core0_ch_outs.v"
`include "dma_axi32_core0_ch_calc.v"
`include "dma_axi32_core0_ch_calc_addr.v"
`include "dma_axi32_core0_ch_calc_size.v"
`include "prgen_min3.v"
`include "prgen_min2.v"
`include "dma_axi32_core0_ch_calc_joint.v"
`include "dma_axi32_core0_ch_periph_mux.v"
`include "dma_axi32_core0_ch_fifo_ctrl.v"
`include "dma_axi32_core0_ch_wr_slicer.v"
`include "prgen_swap_32.v"
`include "dma_axi32_core0_ch_rd_slicer.v"
`include "dma_axi32_core0_ch_fifo_ptr.v"
`include "dma_axi32_core0_ch_fifo.v"
`include "dma_axi32_core0_ch_empty.v"
`include "prgen_delay.v"